module f2_vram(
input wire [7:0] pixel_addr,
input wire [2:0] image_index,
output reg [2:0] pixel_data);

always @(*) begin
	//Get the image index.
	case (image_index)
		3'b000: begin
			case (pixel_addr)
				0	: pixel_data = 3'b111;
				1	: pixel_data = 3'b111;
				2	: pixel_data = 3'b111;
				3	: pixel_data = 3'b111;
				4	: pixel_data = 3'b111;
				5	: pixel_data = 3'b111;
				6	: pixel_data = 3'b111;
				7	: pixel_data = 3'b111;
				8	: pixel_data = 3'b111;
				9	: pixel_data = 3'b111;
				10	: pixel_data = 3'b111;
				11	: pixel_data = 3'b111;
				12	: pixel_data = 3'b111;
				13	: pixel_data = 3'b111;
				14	: pixel_data = 3'b111;
				15	: pixel_data = 3'b111;
				16	: pixel_data = 3'b111;
				17	: pixel_data = 3'b111;
				18	: pixel_data = 3'b111;
				19	: pixel_data = 3'b111;
				20	: pixel_data = 3'b111;
				21	: pixel_data = 3'b111;
				22	: pixel_data = 3'b000;
				23	: pixel_data = 3'b000;
				24	: pixel_data = 3'b000;
				25	: pixel_data = 3'b000;
				26	: pixel_data = 3'b111;
				27	: pixel_data = 3'b111;
				28	: pixel_data = 3'b111;
				29	: pixel_data = 3'b111;
				30	: pixel_data = 3'b111;
				31	: pixel_data = 3'b111;
				32	: pixel_data = 3'b111;
				33	: pixel_data = 3'b111;
				34	: pixel_data = 3'b111;
				35	: pixel_data = 3'b111;
				36	: pixel_data = 3'b111;
				37	: pixel_data = 3'b000;
				38	: pixel_data = 3'b000;
				39	: pixel_data = 3'b000;
				40	: pixel_data = 3'b000;
				41	: pixel_data = 3'b000;
				42	: pixel_data = 3'b000;
				43	: pixel_data = 3'b111;
				44	: pixel_data = 3'b111;
				45	: pixel_data = 3'b111;
				46	: pixel_data = 3'b111;
				47	: pixel_data = 3'b111;
				48	: pixel_data = 3'b111;
				49	: pixel_data = 3'b111;
				50	: pixel_data = 3'b111;
				51	: pixel_data = 3'b111;
				52	: pixel_data = 3'b000;
				53	: pixel_data = 3'b000;
				54	: pixel_data = 3'b111;
				55	: pixel_data = 3'b111;
				56	: pixel_data = 3'b111;
				57	: pixel_data = 3'b111;
				58	: pixel_data = 3'b000;
				59	: pixel_data = 3'b000;
				60	: pixel_data = 3'b111;
				61	: pixel_data = 3'b111;
				62	: pixel_data = 3'b111;
				63	: pixel_data = 3'b111;
				64	: pixel_data = 3'b111;
				65	: pixel_data = 3'b111;
				66	: pixel_data = 3'b111;
				67	: pixel_data = 3'b111;
				68	: pixel_data = 3'b000;
				69	: pixel_data = 3'b111;
				70	: pixel_data = 3'b111;
				71	: pixel_data = 3'b111;
				72	: pixel_data = 3'b111;
				73	: pixel_data = 3'b111;
				74	: pixel_data = 3'b111;
				75	: pixel_data = 3'b000;
				76	: pixel_data = 3'b111;
				77	: pixel_data = 3'b111;
				78	: pixel_data = 3'b111;
				79	: pixel_data = 3'b111;
				80	: pixel_data = 3'b111;
				81	: pixel_data = 3'b111;
				82	: pixel_data = 3'b111;
				83	: pixel_data = 3'b111;
				84	: pixel_data = 3'b000;
				85	: pixel_data = 3'b111;
				86	: pixel_data = 3'b000;
				87	: pixel_data = 3'b111;
				88	: pixel_data = 3'b111;
				89	: pixel_data = 3'b000;
				90	: pixel_data = 3'b111;
				91	: pixel_data = 3'b000;
				92	: pixel_data = 3'b111;
				93	: pixel_data = 3'b111;
				94	: pixel_data = 3'b111;
				95	: pixel_data = 3'b111;
				96	: pixel_data = 3'b111;
				97	: pixel_data = 3'b111;
				98	: pixel_data = 3'b111;
				99	: pixel_data = 3'b000;
				100	: pixel_data = 3'b000;
				101	: pixel_data = 3'b111;
				102	: pixel_data = 3'b000;
				103	: pixel_data = 3'b111;
				104	: pixel_data = 3'b111;
				105	: pixel_data = 3'b000;
				106	: pixel_data = 3'b111;
				107	: pixel_data = 3'b000;
				108	: pixel_data = 3'b000;
				109	: pixel_data = 3'b111;
				110	: pixel_data = 3'b111;
				111	: pixel_data = 3'b111;
				112	: pixel_data = 3'b111;
				113	: pixel_data = 3'b111;
				114	: pixel_data = 3'b000;
				115	: pixel_data = 3'b000;
				116	: pixel_data = 3'b111;
				117	: pixel_data = 3'b111;
				118	: pixel_data = 3'b111;
				119	: pixel_data = 3'b110;
				120	: pixel_data = 3'b110;
				121	: pixel_data = 3'b111;
				122	: pixel_data = 3'b111;
				123	: pixel_data = 3'b111;
				124	: pixel_data = 3'b000;
				125	: pixel_data = 3'b000;
				126	: pixel_data = 3'b111;
				127	: pixel_data = 3'b111;
				128	: pixel_data = 3'b111;
				129	: pixel_data = 3'b111;
				130	: pixel_data = 3'b000;
				131	: pixel_data = 3'b000;
				132	: pixel_data = 3'b111;
				133	: pixel_data = 3'b111;
				134	: pixel_data = 3'b111;
				135	: pixel_data = 3'b111;
				136	: pixel_data = 3'b111;
				137	: pixel_data = 3'b111;
				138	: pixel_data = 3'b111;
				139	: pixel_data = 3'b111;
				140	: pixel_data = 3'b000;
				141	: pixel_data = 3'b000;
				142	: pixel_data = 3'b111;
				143	: pixel_data = 3'b111;
				144	: pixel_data = 3'b111;
				145	: pixel_data = 3'b111;
				146	: pixel_data = 3'b000;
				147	: pixel_data = 3'b000;
				148	: pixel_data = 3'b111;
				149	: pixel_data = 3'b111;
				150	: pixel_data = 3'b111;
				151	: pixel_data = 3'b111;
				152	: pixel_data = 3'b111;
				153	: pixel_data = 3'b111;
				154	: pixel_data = 3'b111;
				155	: pixel_data = 3'b111;
				156	: pixel_data = 3'b000;
				157	: pixel_data = 3'b000;
				158	: pixel_data = 3'b111;
				159	: pixel_data = 3'b111;
				160	: pixel_data = 3'b111;
				161	: pixel_data = 3'b111;
				162	: pixel_data = 3'b111;
				163	: pixel_data = 3'b000;
				164	: pixel_data = 3'b000;
				165	: pixel_data = 3'b111;
				166	: pixel_data = 3'b111;
				167	: pixel_data = 3'b111;
				168	: pixel_data = 3'b111;
				169	: pixel_data = 3'b111;
				170	: pixel_data = 3'b111;
				171	: pixel_data = 3'b000;
				172	: pixel_data = 3'b000;
				173	: pixel_data = 3'b111;
				174	: pixel_data = 3'b111;
				175	: pixel_data = 3'b111;
				176	: pixel_data = 3'b111;
				177	: pixel_data = 3'b111;
				178	: pixel_data = 3'b111;
				179	: pixel_data = 3'b111;
				180	: pixel_data = 3'b000;
				181	: pixel_data = 3'b111;
				182	: pixel_data = 3'b111;
				183	: pixel_data = 3'b111;
				184	: pixel_data = 3'b111;
				185	: pixel_data = 3'b111;
				186	: pixel_data = 3'b111;
				187	: pixel_data = 3'b000;
				188	: pixel_data = 3'b111;
				189	: pixel_data = 3'b111;
				190	: pixel_data = 3'b111;
				191	: pixel_data = 3'b111;
				192	: pixel_data = 3'b111;
				193	: pixel_data = 3'b111;
				194	: pixel_data = 3'b111;
				195	: pixel_data = 3'b111;
				196	: pixel_data = 3'b000;
				197	: pixel_data = 3'b111;
				198	: pixel_data = 3'b111;
				199	: pixel_data = 3'b111;
				200	: pixel_data = 3'b111;
				201	: pixel_data = 3'b111;
				202	: pixel_data = 3'b111;
				203	: pixel_data = 3'b000;
				204	: pixel_data = 3'b111;
				205	: pixel_data = 3'b111;
				206	: pixel_data = 3'b111;
				207	: pixel_data = 3'b111;
				208	: pixel_data = 3'b111;
				209	: pixel_data = 3'b111;
				210	: pixel_data = 3'b111;
				211	: pixel_data = 3'b111;
				212	: pixel_data = 3'b111;
				213	: pixel_data = 3'b110;
				214	: pixel_data = 3'b110;
				215	: pixel_data = 3'b000;
				216	: pixel_data = 3'b000;
				217	: pixel_data = 3'b110;
				218	: pixel_data = 3'b110;
				219	: pixel_data = 3'b111;
				220	: pixel_data = 3'b111;
				221	: pixel_data = 3'b111;
				222	: pixel_data = 3'b111;
				223	: pixel_data = 3'b111;
				224	: pixel_data = 3'b111;
				225	: pixel_data = 3'b111;
				226	: pixel_data = 3'b111;
				227	: pixel_data = 3'b111;
				228	: pixel_data = 3'b111;
				229	: pixel_data = 3'b111;
				230	: pixel_data = 3'b111;
				231	: pixel_data = 3'b111;
				232	: pixel_data = 3'b111;
				233	: pixel_data = 3'b111;
				234	: pixel_data = 3'b111;
				235	: pixel_data = 3'b111;
				236	: pixel_data = 3'b111;
				237	: pixel_data = 3'b111;
				238	: pixel_data = 3'b111;
				239	: pixel_data = 3'b111;
				240	: pixel_data = 3'b111;
				241	: pixel_data = 3'b111;
				242	: pixel_data = 3'b111;
				243	: pixel_data = 3'b111;
				244	: pixel_data = 3'b111;
				245	: pixel_data = 3'b111;
				246	: pixel_data = 3'b111;
				247	: pixel_data = 3'b111;
				248	: pixel_data = 3'b111;
				249	: pixel_data = 3'b111;
				250	: pixel_data = 3'b111;
				251	: pixel_data = 3'b111;
				252	: pixel_data = 3'b111;
				253	: pixel_data = 3'b111;
				254	: pixel_data = 3'b111;
				255	: pixel_data = 3'b111;
			endcase
		end
		3'b001: begin
			case (pixel_addr)
				0	: pixel_data = 3'b111;
				1	: pixel_data = 3'b111;
				2	: pixel_data = 3'b111;
				3	: pixel_data = 3'b111;
				4	: pixel_data = 3'b111;
				5	: pixel_data = 3'b111;
				6	: pixel_data = 3'b111;
				7	: pixel_data = 3'b111;
				8	: pixel_data = 3'b111;
				9	: pixel_data = 3'b111;
				10	: pixel_data = 3'b111;
				11	: pixel_data = 3'b111;
				12	: pixel_data = 3'b111;
				13	: pixel_data = 3'b111;
				14	: pixel_data = 3'b111;
				15	: pixel_data = 3'b111;
				16	: pixel_data = 3'b111;
				17	: pixel_data = 3'b111;
				18	: pixel_data = 3'b111;
				19	: pixel_data = 3'b111;
				20	: pixel_data = 3'b111;
				21	: pixel_data = 3'b111;
				22	: pixel_data = 3'b000;
				23	: pixel_data = 3'b000;
				24	: pixel_data = 3'b000;
				25	: pixel_data = 3'b000;
				26	: pixel_data = 3'b111;
				27	: pixel_data = 3'b111;
				28	: pixel_data = 3'b111;
				29	: pixel_data = 3'b111;
				30	: pixel_data = 3'b111;
				31	: pixel_data = 3'b111;
				32	: pixel_data = 3'b111;
				33	: pixel_data = 3'b111;
				34	: pixel_data = 3'b111;
				35	: pixel_data = 3'b111;
				36	: pixel_data = 3'b111;
				37	: pixel_data = 3'b000;
				38	: pixel_data = 3'b000;
				39	: pixel_data = 3'b000;
				40	: pixel_data = 3'b000;
				41	: pixel_data = 3'b000;
				42	: pixel_data = 3'b000;
				43	: pixel_data = 3'b111;
				44	: pixel_data = 3'b111;
				45	: pixel_data = 3'b111;
				46	: pixel_data = 3'b111;
				47	: pixel_data = 3'b111;
				48	: pixel_data = 3'b111;
				49	: pixel_data = 3'b111;
				50	: pixel_data = 3'b111;
				51	: pixel_data = 3'b111;
				52	: pixel_data = 3'b111;
				53	: pixel_data = 3'b000;
				54	: pixel_data = 3'b111;
				55	: pixel_data = 3'b111;
				56	: pixel_data = 3'b111;
				57	: pixel_data = 3'b111;
				58	: pixel_data = 3'b000;
				59	: pixel_data = 3'b111;
				60	: pixel_data = 3'b111;
				61	: pixel_data = 3'b111;
				62	: pixel_data = 3'b111;
				63	: pixel_data = 3'b111;
				64	: pixel_data = 3'b111;
				65	: pixel_data = 3'b111;
				66	: pixel_data = 3'b111;
				67	: pixel_data = 3'b111;
				68	: pixel_data = 3'b111;
				69	: pixel_data = 3'b000;
				70	: pixel_data = 3'b111;
				71	: pixel_data = 3'b000;
				72	: pixel_data = 3'b111;
				73	: pixel_data = 3'b111;
				74	: pixel_data = 3'b000;
				75	: pixel_data = 3'b111;
				76	: pixel_data = 3'b111;
				77	: pixel_data = 3'b111;
				78	: pixel_data = 3'b111;
				79	: pixel_data = 3'b111;
				80	: pixel_data = 3'b111;
				81	: pixel_data = 3'b111;
				82	: pixel_data = 3'b111;
				83	: pixel_data = 3'b111;
				84	: pixel_data = 3'b111;
				85	: pixel_data = 3'b000;
				86	: pixel_data = 3'b111;
				87	: pixel_data = 3'b000;
				88	: pixel_data = 3'b111;
				89	: pixel_data = 3'b111;
				90	: pixel_data = 3'b000;
				91	: pixel_data = 3'b111;
				92	: pixel_data = 3'b111;
				93	: pixel_data = 3'b111;
				94	: pixel_data = 3'b111;
				95	: pixel_data = 3'b111;
				96	: pixel_data = 3'b111;
				97	: pixel_data = 3'b111;
				98	: pixel_data = 3'b111;
				99	: pixel_data = 3'b111;
				100	: pixel_data = 3'b110;
				101	: pixel_data = 3'b110;
				102	: pixel_data = 3'b111;
				103	: pixel_data = 3'b111;
				104	: pixel_data = 3'b111;
				105	: pixel_data = 3'b111;
				106	: pixel_data = 3'b000;
				107	: pixel_data = 3'b111;
				108	: pixel_data = 3'b111;
				109	: pixel_data = 3'b111;
				110	: pixel_data = 3'b111;
				111	: pixel_data = 3'b111;
				112	: pixel_data = 3'b111;
				113	: pixel_data = 3'b111;
				114	: pixel_data = 3'b111;
				115	: pixel_data = 3'b111;
				116	: pixel_data = 3'b111;
				117	: pixel_data = 3'b000;
				118	: pixel_data = 3'b111;
				119	: pixel_data = 3'b000;
				120	: pixel_data = 3'b000;
				121	: pixel_data = 3'b000;
				122	: pixel_data = 3'b000;
				123	: pixel_data = 3'b111;
				124	: pixel_data = 3'b111;
				125	: pixel_data = 3'b111;
				126	: pixel_data = 3'b111;
				127	: pixel_data = 3'b111;
				128	: pixel_data = 3'b111;
				129	: pixel_data = 3'b111;
				130	: pixel_data = 3'b111;
				131	: pixel_data = 3'b111;
				132	: pixel_data = 3'b111;
				133	: pixel_data = 3'b000;
				134	: pixel_data = 3'b111;
				135	: pixel_data = 3'b000;
				136	: pixel_data = 3'b000;
				137	: pixel_data = 3'b000;
				138	: pixel_data = 3'b111;
				139	: pixel_data = 3'b111;
				140	: pixel_data = 3'b111;
				141	: pixel_data = 3'b111;
				142	: pixel_data = 3'b111;
				143	: pixel_data = 3'b111;
				144	: pixel_data = 3'b111;
				145	: pixel_data = 3'b111;
				146	: pixel_data = 3'b111;
				147	: pixel_data = 3'b111;
				148	: pixel_data = 3'b111;
				149	: pixel_data = 3'b000;
				150	: pixel_data = 3'b111;
				151	: pixel_data = 3'b000;
				152	: pixel_data = 3'b000;
				153	: pixel_data = 3'b000;
				154	: pixel_data = 3'b111;
				155	: pixel_data = 3'b111;
				156	: pixel_data = 3'b111;
				157	: pixel_data = 3'b111;
				158	: pixel_data = 3'b111;
				159	: pixel_data = 3'b111;
				160	: pixel_data = 3'b111;
				161	: pixel_data = 3'b111;
				162	: pixel_data = 3'b111;
				163	: pixel_data = 3'b111;
				164	: pixel_data = 3'b111;
				165	: pixel_data = 3'b000;
				166	: pixel_data = 3'b111;
				167	: pixel_data = 3'b000;
				168	: pixel_data = 3'b111;
				169	: pixel_data = 3'b000;
				170	: pixel_data = 3'b111;
				171	: pixel_data = 3'b111;
				172	: pixel_data = 3'b111;
				173	: pixel_data = 3'b111;
				174	: pixel_data = 3'b111;
				175	: pixel_data = 3'b111;
				176	: pixel_data = 3'b111;
				177	: pixel_data = 3'b111;
				178	: pixel_data = 3'b111;
				179	: pixel_data = 3'b111;
				180	: pixel_data = 3'b111;
				181	: pixel_data = 3'b000;
				182	: pixel_data = 3'b111;
				183	: pixel_data = 3'b111;
				184	: pixel_data = 3'b111;
				185	: pixel_data = 3'b000;
				186	: pixel_data = 3'b111;
				187	: pixel_data = 3'b111;
				188	: pixel_data = 3'b111;
				189	: pixel_data = 3'b111;
				190	: pixel_data = 3'b111;
				191	: pixel_data = 3'b111;
				192	: pixel_data = 3'b111;
				193	: pixel_data = 3'b111;
				194	: pixel_data = 3'b111;
				195	: pixel_data = 3'b111;
				196	: pixel_data = 3'b111;
				197	: pixel_data = 3'b000;
				198	: pixel_data = 3'b111;
				199	: pixel_data = 3'b111;
				200	: pixel_data = 3'b000;
				201	: pixel_data = 3'b000;
				202	: pixel_data = 3'b111;
				203	: pixel_data = 3'b111;
				204	: pixel_data = 3'b111;
				205	: pixel_data = 3'b111;
				206	: pixel_data = 3'b111;
				207	: pixel_data = 3'b111;
				208	: pixel_data = 3'b111;
				209	: pixel_data = 3'b111;
				210	: pixel_data = 3'b111;
				211	: pixel_data = 3'b111;
				212	: pixel_data = 3'b110;
				213	: pixel_data = 3'b110;
				214	: pixel_data = 3'b000;
				215	: pixel_data = 3'b000;
				216	: pixel_data = 3'b000;
				217	: pixel_data = 3'b111;
				218	: pixel_data = 3'b111;
				219	: pixel_data = 3'b111;
				220	: pixel_data = 3'b111;
				221	: pixel_data = 3'b111;
				222	: pixel_data = 3'b111;
				223	: pixel_data = 3'b111;
				224	: pixel_data = 3'b111;
				225	: pixel_data = 3'b111;
				226	: pixel_data = 3'b111;
				227	: pixel_data = 3'b111;
				228	: pixel_data = 3'b111;
				229	: pixel_data = 3'b111;
				230	: pixel_data = 3'b111;
				231	: pixel_data = 3'b111;
				232	: pixel_data = 3'b111;
				233	: pixel_data = 3'b111;
				234	: pixel_data = 3'b111;
				235	: pixel_data = 3'b111;
				236	: pixel_data = 3'b111;
				237	: pixel_data = 3'b111;
				238	: pixel_data = 3'b111;
				239	: pixel_data = 3'b111;
				240	: pixel_data = 3'b111;
				241	: pixel_data = 3'b111;
				242	: pixel_data = 3'b111;
				243	: pixel_data = 3'b111;
				244	: pixel_data = 3'b111;
				245	: pixel_data = 3'b111;
				246	: pixel_data = 3'b111;
				247	: pixel_data = 3'b111;
				248	: pixel_data = 3'b111;
				249	: pixel_data = 3'b111;
				250	: pixel_data = 3'b111;
				251	: pixel_data = 3'b111;
				252	: pixel_data = 3'b111;
				253	: pixel_data = 3'b111;
				254	: pixel_data = 3'b111;
				255	: pixel_data = 3'b111;
			endcase
		end
	endcase
end

endmodule