module img_vrom(
input wire [7:0] func2_pixel_addr,
input wire [7:0] func3_pixel_addr,
input wire [2:0] image_index,
output reg [2:0] func2_pixel_data,
output reg [2:0] func3_pixel_data);

reg [2:0] current_image;
reg am, bm, cm;
reg[1:0] dm;

task image0_data;
	input [7:0] image_pixel_addr;
	output [2:0] image_pixel_data;
	reg [2:0] image_pixel_data;
	begin
		case (image_pixel_addr)
			0	: image_pixel_data = 3'b111;
			1	: image_pixel_data = 3'b111;
			2	: image_pixel_data = 3'b111;
			3	: image_pixel_data = 3'b111;
			4	: image_pixel_data = 3'b111;
			5	: image_pixel_data = 3'b111;
			6	: image_pixel_data = 3'b111;
			7	: image_pixel_data = 3'b111;
			8	: image_pixel_data = 3'b111;
			9	: image_pixel_data = 3'b111;
			10	: image_pixel_data = 3'b111;
			11	: image_pixel_data = 3'b111;
			12	: image_pixel_data = 3'b111;
			13	: image_pixel_data = 3'b111;
			14	: image_pixel_data = 3'b111;
			15	: image_pixel_data = 3'b111;
			16	: image_pixel_data = 3'b111;
			17	: image_pixel_data = 3'b111;
			18	: image_pixel_data = 3'b111;
			19	: image_pixel_data = 3'b111;
			20	: image_pixel_data = 3'b111;
			21	: image_pixel_data = 3'b111;
			22	: image_pixel_data = 3'b000;
			23	: image_pixel_data = 3'b000;
			24	: image_pixel_data = 3'b000;
			25	: image_pixel_data = 3'b000;
			26	: image_pixel_data = 3'b111;
			27	: image_pixel_data = 3'b111;
			28	: image_pixel_data = 3'b111;
			29	: image_pixel_data = 3'b111;
			30	: image_pixel_data = 3'b111;
			31	: image_pixel_data = 3'b111;
			32	: image_pixel_data = 3'b111;
			33	: image_pixel_data = 3'b111;
			34	: image_pixel_data = 3'b111;
			35	: image_pixel_data = 3'b111;
			36	: image_pixel_data = 3'b111;
			37	: image_pixel_data = 3'b000;
			38	: image_pixel_data = 3'b000;
			39	: image_pixel_data = 3'b000;
			40	: image_pixel_data = 3'b000;
			41	: image_pixel_data = 3'b000;
			42	: image_pixel_data = 3'b000;
			43	: image_pixel_data = 3'b111;
			44	: image_pixel_data = 3'b111;
			45	: image_pixel_data = 3'b111;
			46	: image_pixel_data = 3'b111;
			47	: image_pixel_data = 3'b111;
			48	: image_pixel_data = 3'b111;
			49	: image_pixel_data = 3'b111;
			50	: image_pixel_data = 3'b111;
			51	: image_pixel_data = 3'b111;
			52	: image_pixel_data = 3'b000;
			53	: image_pixel_data = 3'b000;
			54	: image_pixel_data = 3'b111;
			55	: image_pixel_data = 3'b111;
			56	: image_pixel_data = 3'b111;
			57	: image_pixel_data = 3'b111;
			58	: image_pixel_data = 3'b000;
			59	: image_pixel_data = 3'b000;
			60	: image_pixel_data = 3'b111;
			61	: image_pixel_data = 3'b111;
			62	: image_pixel_data = 3'b111;
			63	: image_pixel_data = 3'b111;
			64	: image_pixel_data = 3'b111;
			65	: image_pixel_data = 3'b111;
			66	: image_pixel_data = 3'b111;
			67	: image_pixel_data = 3'b111;
			68	: image_pixel_data = 3'b000;
			69	: image_pixel_data = 3'b111;
			70	: image_pixel_data = 3'b111;
			71	: image_pixel_data = 3'b111;
			72	: image_pixel_data = 3'b111;
			73	: image_pixel_data = 3'b111;
			74	: image_pixel_data = 3'b111;
			75	: image_pixel_data = 3'b000;
			76	: image_pixel_data = 3'b111;
			77	: image_pixel_data = 3'b111;
			78	: image_pixel_data = 3'b111;
			79	: image_pixel_data = 3'b111;
			80	: image_pixel_data = 3'b111;
			81	: image_pixel_data = 3'b111;
			82	: image_pixel_data = 3'b111;
			83	: image_pixel_data = 3'b111;
			84	: image_pixel_data = 3'b000;
			85	: image_pixel_data = 3'b111;
			86	: image_pixel_data = 3'b000;
			87	: image_pixel_data = 3'b111;
			88	: image_pixel_data = 3'b111;
			89	: image_pixel_data = 3'b000;
			90	: image_pixel_data = 3'b111;
			91	: image_pixel_data = 3'b000;
			92	: image_pixel_data = 3'b111;
			93	: image_pixel_data = 3'b111;
			94	: image_pixel_data = 3'b111;
			95	: image_pixel_data = 3'b111;
			96	: image_pixel_data = 3'b111;
			97	: image_pixel_data = 3'b111;
			98	: image_pixel_data = 3'b111;
			99	: image_pixel_data = 3'b000;
			100	: image_pixel_data = 3'b000;
			101	: image_pixel_data = 3'b111;
			102	: image_pixel_data = 3'b000;
			103	: image_pixel_data = 3'b111;
			104	: image_pixel_data = 3'b111;
			105	: image_pixel_data = 3'b000;
			106	: image_pixel_data = 3'b111;
			107	: image_pixel_data = 3'b000;
			108	: image_pixel_data = 3'b000;
			109	: image_pixel_data = 3'b111;
			110	: image_pixel_data = 3'b111;
			111	: image_pixel_data = 3'b111;
			112	: image_pixel_data = 3'b111;
			113	: image_pixel_data = 3'b111;
			114	: image_pixel_data = 3'b000;
			115	: image_pixel_data = 3'b000;
			116	: image_pixel_data = 3'b111;
			117	: image_pixel_data = 3'b111;
			118	: image_pixel_data = 3'b111;
			119	: image_pixel_data = 3'b110;
			120	: image_pixel_data = 3'b110;
			121	: image_pixel_data = 3'b111;
			122	: image_pixel_data = 3'b111;
			123	: image_pixel_data = 3'b111;
			124	: image_pixel_data = 3'b000;
			125	: image_pixel_data = 3'b000;
			126	: image_pixel_data = 3'b111;
			127	: image_pixel_data = 3'b111;
			128	: image_pixel_data = 3'b111;
			129	: image_pixel_data = 3'b111;
			130	: image_pixel_data = 3'b000;
			131	: image_pixel_data = 3'b000;
			132	: image_pixel_data = 3'b111;
			133	: image_pixel_data = 3'b111;
			134	: image_pixel_data = 3'b111;
			135	: image_pixel_data = 3'b111;
			136	: image_pixel_data = 3'b111;
			137	: image_pixel_data = 3'b111;
			138	: image_pixel_data = 3'b111;
			139	: image_pixel_data = 3'b111;
			140	: image_pixel_data = 3'b000;
			141	: image_pixel_data = 3'b000;
			142	: image_pixel_data = 3'b111;
			143	: image_pixel_data = 3'b111;
			144	: image_pixel_data = 3'b111;
			145	: image_pixel_data = 3'b111;
			146	: image_pixel_data = 3'b000;
			147	: image_pixel_data = 3'b000;
			148	: image_pixel_data = 3'b111;
			149	: image_pixel_data = 3'b111;
			150	: image_pixel_data = 3'b111;
			151	: image_pixel_data = 3'b111;
			152	: image_pixel_data = 3'b111;
			153	: image_pixel_data = 3'b111;
			154	: image_pixel_data = 3'b111;
			155	: image_pixel_data = 3'b111;
			156	: image_pixel_data = 3'b000;
			157	: image_pixel_data = 3'b000;
			158	: image_pixel_data = 3'b111;
			159	: image_pixel_data = 3'b111;
			160	: image_pixel_data = 3'b111;
			161	: image_pixel_data = 3'b111;
			162	: image_pixel_data = 3'b111;
			163	: image_pixel_data = 3'b000;
			164	: image_pixel_data = 3'b000;
			165	: image_pixel_data = 3'b111;
			166	: image_pixel_data = 3'b111;
			167	: image_pixel_data = 3'b111;
			168	: image_pixel_data = 3'b111;
			169	: image_pixel_data = 3'b111;
			170	: image_pixel_data = 3'b111;
			171	: image_pixel_data = 3'b000;
			172	: image_pixel_data = 3'b000;
			173	: image_pixel_data = 3'b111;
			174	: image_pixel_data = 3'b111;
			175	: image_pixel_data = 3'b111;
			176	: image_pixel_data = 3'b111;
			177	: image_pixel_data = 3'b111;
			178	: image_pixel_data = 3'b111;
			179	: image_pixel_data = 3'b111;
			180	: image_pixel_data = 3'b000;
			181	: image_pixel_data = 3'b111;
			182	: image_pixel_data = 3'b111;
			183	: image_pixel_data = 3'b111;
			184	: image_pixel_data = 3'b111;
			185	: image_pixel_data = 3'b111;
			186	: image_pixel_data = 3'b111;
			187	: image_pixel_data = 3'b000;
			188	: image_pixel_data = 3'b111;
			189	: image_pixel_data = 3'b111;
			190	: image_pixel_data = 3'b111;
			191	: image_pixel_data = 3'b111;
			192	: image_pixel_data = 3'b111;
			193	: image_pixel_data = 3'b111;
			194	: image_pixel_data = 3'b111;
			195	: image_pixel_data = 3'b111;
			196	: image_pixel_data = 3'b000;
			197	: image_pixel_data = 3'b111;
			198	: image_pixel_data = 3'b111;
			199	: image_pixel_data = 3'b111;
			200	: image_pixel_data = 3'b111;
			201	: image_pixel_data = 3'b111;
			202	: image_pixel_data = 3'b111;
			203	: image_pixel_data = 3'b000;
			204	: image_pixel_data = 3'b111;
			205	: image_pixel_data = 3'b111;
			206	: image_pixel_data = 3'b111;
			207	: image_pixel_data = 3'b111;
			208	: image_pixel_data = 3'b111;
			209	: image_pixel_data = 3'b111;
			210	: image_pixel_data = 3'b111;
			211	: image_pixel_data = 3'b111;
			212	: image_pixel_data = 3'b111;
			213	: image_pixel_data = 3'b110;
			214	: image_pixel_data = 3'b110;
			215	: image_pixel_data = 3'b000;
			216	: image_pixel_data = 3'b000;
			217	: image_pixel_data = 3'b110;
			218	: image_pixel_data = 3'b110;
			219	: image_pixel_data = 3'b111;
			220	: image_pixel_data = 3'b111;
			221	: image_pixel_data = 3'b111;
			222	: image_pixel_data = 3'b111;
			223	: image_pixel_data = 3'b111;
			224	: image_pixel_data = 3'b111;
			225	: image_pixel_data = 3'b111;
			226	: image_pixel_data = 3'b111;
			227	: image_pixel_data = 3'b111;
			228	: image_pixel_data = 3'b111;
			229	: image_pixel_data = 3'b111;
			230	: image_pixel_data = 3'b111;
			231	: image_pixel_data = 3'b111;
			232	: image_pixel_data = 3'b111;
			233	: image_pixel_data = 3'b111;
			234	: image_pixel_data = 3'b111;
			235	: image_pixel_data = 3'b111;
			236	: image_pixel_data = 3'b111;
			237	: image_pixel_data = 3'b111;
			238	: image_pixel_data = 3'b111;
			239	: image_pixel_data = 3'b111;
			240	: image_pixel_data = 3'b111;
			241	: image_pixel_data = 3'b111;
			242	: image_pixel_data = 3'b111;
			243	: image_pixel_data = 3'b111;
			244	: image_pixel_data = 3'b111;
			245	: image_pixel_data = 3'b111;
			246	: image_pixel_data = 3'b111;
			247	: image_pixel_data = 3'b111;
			248	: image_pixel_data = 3'b111;
			249	: image_pixel_data = 3'b111;
			250	: image_pixel_data = 3'b111;
			251	: image_pixel_data = 3'b111;
			252	: image_pixel_data = 3'b111;
			253	: image_pixel_data = 3'b111;
			254	: image_pixel_data = 3'b111;
			255	: image_pixel_data = 3'b111;
		endcase
	end
endtask

task image1_data;
	input [7:0] image_pixel_addr;
	output [2:0] image_pixel_data;
	reg [2:0] image_pixel_data;
	begin
		case (image_pixel_addr)
			0	: image_pixel_data = 3'b111;
			1	: image_pixel_data = 3'b111;
			2	: image_pixel_data = 3'b111;
			3	: image_pixel_data = 3'b111;
			4	: image_pixel_data = 3'b111;
			5	: image_pixel_data = 3'b111;
			6	: image_pixel_data = 3'b111;
			7	: image_pixel_data = 3'b111;
			8	: image_pixel_data = 3'b111;
			9	: image_pixel_data = 3'b111;
			10	: image_pixel_data = 3'b111;
			11	: image_pixel_data = 3'b111;
			12	: image_pixel_data = 3'b111;
			13	: image_pixel_data = 3'b111;
			14	: image_pixel_data = 3'b111;
			15	: image_pixel_data = 3'b111;
			16	: image_pixel_data = 3'b111;
			17	: image_pixel_data = 3'b111;
			18	: image_pixel_data = 3'b111;
			19	: image_pixel_data = 3'b111;
			20	: image_pixel_data = 3'b111;
			21	: image_pixel_data = 3'b111;
			22	: image_pixel_data = 3'b000;
			23	: image_pixel_data = 3'b000;
			24	: image_pixel_data = 3'b000;
			25	: image_pixel_data = 3'b000;
			26	: image_pixel_data = 3'b111;
			27	: image_pixel_data = 3'b111;
			28	: image_pixel_data = 3'b111;
			29	: image_pixel_data = 3'b111;
			30	: image_pixel_data = 3'b111;
			31	: image_pixel_data = 3'b111;
			32	: image_pixel_data = 3'b111;
			33	: image_pixel_data = 3'b111;
			34	: image_pixel_data = 3'b111;
			35	: image_pixel_data = 3'b111;
			36	: image_pixel_data = 3'b111;
			37	: image_pixel_data = 3'b000;
			38	: image_pixel_data = 3'b000;
			39	: image_pixel_data = 3'b000;
			40	: image_pixel_data = 3'b000;
			41	: image_pixel_data = 3'b000;
			42	: image_pixel_data = 3'b000;
			43	: image_pixel_data = 3'b111;
			44	: image_pixel_data = 3'b111;
			45	: image_pixel_data = 3'b111;
			46	: image_pixel_data = 3'b111;
			47	: image_pixel_data = 3'b111;
			48	: image_pixel_data = 3'b111;
			49	: image_pixel_data = 3'b111;
			50	: image_pixel_data = 3'b111;
			51	: image_pixel_data = 3'b111;
			52	: image_pixel_data = 3'b111;
			53	: image_pixel_data = 3'b000;
			54	: image_pixel_data = 3'b111;
			55	: image_pixel_data = 3'b111;
			56	: image_pixel_data = 3'b111;
			57	: image_pixel_data = 3'b111;
			58	: image_pixel_data = 3'b000;
			59	: image_pixel_data = 3'b111;
			60	: image_pixel_data = 3'b111;
			61	: image_pixel_data = 3'b111;
			62	: image_pixel_data = 3'b111;
			63	: image_pixel_data = 3'b111;
			64	: image_pixel_data = 3'b111;
			65	: image_pixel_data = 3'b111;
			66	: image_pixel_data = 3'b111;
			67	: image_pixel_data = 3'b111;
			68	: image_pixel_data = 3'b111;
			69	: image_pixel_data = 3'b000;
			70	: image_pixel_data = 3'b111;
			71	: image_pixel_data = 3'b000;
			72	: image_pixel_data = 3'b111;
			73	: image_pixel_data = 3'b111;
			74	: image_pixel_data = 3'b000;
			75	: image_pixel_data = 3'b111;
			76	: image_pixel_data = 3'b111;
			77	: image_pixel_data = 3'b111;
			78	: image_pixel_data = 3'b111;
			79	: image_pixel_data = 3'b111;
			80	: image_pixel_data = 3'b111;
			81	: image_pixel_data = 3'b111;
			82	: image_pixel_data = 3'b111;
			83	: image_pixel_data = 3'b111;
			84	: image_pixel_data = 3'b111;
			85	: image_pixel_data = 3'b000;
			86	: image_pixel_data = 3'b111;
			87	: image_pixel_data = 3'b000;
			88	: image_pixel_data = 3'b111;
			89	: image_pixel_data = 3'b111;
			90	: image_pixel_data = 3'b000;
			91	: image_pixel_data = 3'b111;
			92	: image_pixel_data = 3'b111;
			93	: image_pixel_data = 3'b111;
			94	: image_pixel_data = 3'b111;
			95	: image_pixel_data = 3'b111;
			96	: image_pixel_data = 3'b111;
			97	: image_pixel_data = 3'b111;
			98	: image_pixel_data = 3'b111;
			99	: image_pixel_data = 3'b111;
			100	: image_pixel_data = 3'b110;
			101	: image_pixel_data = 3'b110;
			102	: image_pixel_data = 3'b111;
			103	: image_pixel_data = 3'b111;
			104	: image_pixel_data = 3'b111;
			105	: image_pixel_data = 3'b111;
			106	: image_pixel_data = 3'b000;
			107	: image_pixel_data = 3'b111;
			108	: image_pixel_data = 3'b111;
			109	: image_pixel_data = 3'b111;
			110	: image_pixel_data = 3'b111;
			111	: image_pixel_data = 3'b111;
			112	: image_pixel_data = 3'b111;
			113	: image_pixel_data = 3'b111;
			114	: image_pixel_data = 3'b111;
			115	: image_pixel_data = 3'b111;
			116	: image_pixel_data = 3'b111;
			117	: image_pixel_data = 3'b000;
			118	: image_pixel_data = 3'b111;
			119	: image_pixel_data = 3'b000;
			120	: image_pixel_data = 3'b000;
			121	: image_pixel_data = 3'b000;
			122	: image_pixel_data = 3'b000;
			123	: image_pixel_data = 3'b111;
			124	: image_pixel_data = 3'b111;
			125	: image_pixel_data = 3'b111;
			126	: image_pixel_data = 3'b111;
			127	: image_pixel_data = 3'b111;
			128	: image_pixel_data = 3'b111;
			129	: image_pixel_data = 3'b111;
			130	: image_pixel_data = 3'b111;
			131	: image_pixel_data = 3'b111;
			132	: image_pixel_data = 3'b111;
			133	: image_pixel_data = 3'b000;
			134	: image_pixel_data = 3'b111;
			135	: image_pixel_data = 3'b000;
			136	: image_pixel_data = 3'b000;
			137	: image_pixel_data = 3'b000;
			138	: image_pixel_data = 3'b111;
			139	: image_pixel_data = 3'b111;
			140	: image_pixel_data = 3'b111;
			141	: image_pixel_data = 3'b111;
			142	: image_pixel_data = 3'b111;
			143	: image_pixel_data = 3'b111;
			144	: image_pixel_data = 3'b111;
			145	: image_pixel_data = 3'b111;
			146	: image_pixel_data = 3'b111;
			147	: image_pixel_data = 3'b111;
			148	: image_pixel_data = 3'b111;
			149	: image_pixel_data = 3'b000;
			150	: image_pixel_data = 3'b111;
			151	: image_pixel_data = 3'b000;
			152	: image_pixel_data = 3'b000;
			153	: image_pixel_data = 3'b000;
			154	: image_pixel_data = 3'b111;
			155	: image_pixel_data = 3'b111;
			156	: image_pixel_data = 3'b111;
			157	: image_pixel_data = 3'b111;
			158	: image_pixel_data = 3'b111;
			159	: image_pixel_data = 3'b111;
			160	: image_pixel_data = 3'b111;
			161	: image_pixel_data = 3'b111;
			162	: image_pixel_data = 3'b111;
			163	: image_pixel_data = 3'b111;
			164	: image_pixel_data = 3'b111;
			165	: image_pixel_data = 3'b000;
			166	: image_pixel_data = 3'b111;
			167	: image_pixel_data = 3'b000;
			168	: image_pixel_data = 3'b111;
			169	: image_pixel_data = 3'b000;
			170	: image_pixel_data = 3'b111;
			171	: image_pixel_data = 3'b111;
			172	: image_pixel_data = 3'b111;
			173	: image_pixel_data = 3'b111;
			174	: image_pixel_data = 3'b111;
			175	: image_pixel_data = 3'b111;
			176	: image_pixel_data = 3'b111;
			177	: image_pixel_data = 3'b111;
			178	: image_pixel_data = 3'b111;
			179	: image_pixel_data = 3'b111;
			180	: image_pixel_data = 3'b111;
			181	: image_pixel_data = 3'b000;
			182	: image_pixel_data = 3'b111;
			183	: image_pixel_data = 3'b111;
			184	: image_pixel_data = 3'b111;
			185	: image_pixel_data = 3'b000;
			186	: image_pixel_data = 3'b111;
			187	: image_pixel_data = 3'b111;
			188	: image_pixel_data = 3'b111;
			189	: image_pixel_data = 3'b111;
			190	: image_pixel_data = 3'b111;
			191	: image_pixel_data = 3'b111;
			192	: image_pixel_data = 3'b111;
			193	: image_pixel_data = 3'b111;
			194	: image_pixel_data = 3'b111;
			195	: image_pixel_data = 3'b111;
			196	: image_pixel_data = 3'b111;
			197	: image_pixel_data = 3'b000;
			198	: image_pixel_data = 3'b111;
			199	: image_pixel_data = 3'b111;
			200	: image_pixel_data = 3'b000;
			201	: image_pixel_data = 3'b000;
			202	: image_pixel_data = 3'b111;
			203	: image_pixel_data = 3'b111;
			204	: image_pixel_data = 3'b111;
			205	: image_pixel_data = 3'b111;
			206	: image_pixel_data = 3'b111;
			207	: image_pixel_data = 3'b111;
			208	: image_pixel_data = 3'b111;
			209	: image_pixel_data = 3'b111;
			210	: image_pixel_data = 3'b111;
			211	: image_pixel_data = 3'b111;
			212	: image_pixel_data = 3'b110;
			213	: image_pixel_data = 3'b110;
			214	: image_pixel_data = 3'b000;
			215	: image_pixel_data = 3'b000;
			216	: image_pixel_data = 3'b000;
			217	: image_pixel_data = 3'b111;
			218	: image_pixel_data = 3'b111;
			219	: image_pixel_data = 3'b111;
			220	: image_pixel_data = 3'b111;
			221	: image_pixel_data = 3'b111;
			222	: image_pixel_data = 3'b111;
			223	: image_pixel_data = 3'b111;
			224	: image_pixel_data = 3'b111;
			225	: image_pixel_data = 3'b111;
			226	: image_pixel_data = 3'b111;
			227	: image_pixel_data = 3'b111;
			228	: image_pixel_data = 3'b111;
			229	: image_pixel_data = 3'b111;
			230	: image_pixel_data = 3'b111;
			231	: image_pixel_data = 3'b111;
			232	: image_pixel_data = 3'b111;
			233	: image_pixel_data = 3'b111;
			234	: image_pixel_data = 3'b111;
			235	: image_pixel_data = 3'b111;
			236	: image_pixel_data = 3'b111;
			237	: image_pixel_data = 3'b111;
			238	: image_pixel_data = 3'b111;
			239	: image_pixel_data = 3'b111;
			240	: image_pixel_data = 3'b111;
			241	: image_pixel_data = 3'b111;
			242	: image_pixel_data = 3'b111;
			243	: image_pixel_data = 3'b111;
			244	: image_pixel_data = 3'b111;
			245	: image_pixel_data = 3'b111;
			246	: image_pixel_data = 3'b111;
			247	: image_pixel_data = 3'b111;
			248	: image_pixel_data = 3'b111;
			249	: image_pixel_data = 3'b111;
			250	: image_pixel_data = 3'b111;
			251	: image_pixel_data = 3'b111;
			252	: image_pixel_data = 3'b111;
			253	: image_pixel_data = 3'b111;
			254	: image_pixel_data = 3'b111;
			255	: image_pixel_data = 3'b111;
		endcase
	end
endtask

task image2_data;
	input [7:0] image_pixel_addr;
	output [2:0] image_pixel_data;
	reg [2:0] image_pixel_data;
	begin
		case (image_pixel_addr)
			0	: image_pixel_data = 3'b111;
			1	: image_pixel_data = 3'b111;
			2	: image_pixel_data = 3'b111;
			3	: image_pixel_data = 3'b111;
			4	: image_pixel_data = 3'b111;
			5	: image_pixel_data = 3'b111;
			6	: image_pixel_data = 3'b111;
			7	: image_pixel_data = 3'b111;
			8	: image_pixel_data = 3'b111;
			9	: image_pixel_data = 3'b111;
			10	: image_pixel_data = 3'b111;
			11	: image_pixel_data = 3'b111;
			12	: image_pixel_data = 3'b111;
			13	: image_pixel_data = 3'b111;
			14	: image_pixel_data = 3'b111;
			15	: image_pixel_data = 3'b111;
			16	: image_pixel_data = 3'b111;
			17	: image_pixel_data = 3'b111;
			18	: image_pixel_data = 3'b111;
			19	: image_pixel_data = 3'b111;
			20	: image_pixel_data = 3'b111;
			21	: image_pixel_data = 3'b111;
			22	: image_pixel_data = 3'b000;
			23	: image_pixel_data = 3'b000;
			24	: image_pixel_data = 3'b000;
			25	: image_pixel_data = 3'b000;
			26	: image_pixel_data = 3'b111;
			27	: image_pixel_data = 3'b111;
			28	: image_pixel_data = 3'b111;
			29	: image_pixel_data = 3'b111;
			30	: image_pixel_data = 3'b111;
			31	: image_pixel_data = 3'b111;
			32	: image_pixel_data = 3'b111;
			33	: image_pixel_data = 3'b111;
			34	: image_pixel_data = 3'b111;
			35	: image_pixel_data = 3'b111;
			36	: image_pixel_data = 3'b111;
			37	: image_pixel_data = 3'b000;
			38	: image_pixel_data = 3'b000;
			39	: image_pixel_data = 3'b111;
			40	: image_pixel_data = 3'b111;
			41	: image_pixel_data = 3'b000;
			42	: image_pixel_data = 3'b000;
			43	: image_pixel_data = 3'b111;
			44	: image_pixel_data = 3'b111;
			45	: image_pixel_data = 3'b111;
			46	: image_pixel_data = 3'b111;
			47	: image_pixel_data = 3'b111;
			48	: image_pixel_data = 3'b111;
			49	: image_pixel_data = 3'b111;
			50	: image_pixel_data = 3'b111;
			51	: image_pixel_data = 3'b111;
			52	: image_pixel_data = 3'b111;
			53	: image_pixel_data = 3'b000;
			54	: image_pixel_data = 3'b111;
			55	: image_pixel_data = 3'b111;
			56	: image_pixel_data = 3'b111;
			57	: image_pixel_data = 3'b111;
			58	: image_pixel_data = 3'b000;
			59	: image_pixel_data = 3'b111;
			60	: image_pixel_data = 3'b111;
			61	: image_pixel_data = 3'b111;
			62	: image_pixel_data = 3'b111;
			63	: image_pixel_data = 3'b111;
			64	: image_pixel_data = 3'b111;
			65	: image_pixel_data = 3'b111;
			66	: image_pixel_data = 3'b111;
			67	: image_pixel_data = 3'b111;
			68	: image_pixel_data = 3'b111;
			69	: image_pixel_data = 3'b000;
			70	: image_pixel_data = 3'b111;
			71	: image_pixel_data = 3'b111;
			72	: image_pixel_data = 3'b000;
			73	: image_pixel_data = 3'b111;
			74	: image_pixel_data = 3'b000;
			75	: image_pixel_data = 3'b111;
			76	: image_pixel_data = 3'b111;
			77	: image_pixel_data = 3'b111;
			78	: image_pixel_data = 3'b111;
			79	: image_pixel_data = 3'b111;
			80	: image_pixel_data = 3'b111;
			81	: image_pixel_data = 3'b111;
			82	: image_pixel_data = 3'b111;
			83	: image_pixel_data = 3'b111;
			84	: image_pixel_data = 3'b111;
			85	: image_pixel_data = 3'b000;
			86	: image_pixel_data = 3'b111;
			87	: image_pixel_data = 3'b111;
			88	: image_pixel_data = 3'b000;
			89	: image_pixel_data = 3'b111;
			90	: image_pixel_data = 3'b000;
			91	: image_pixel_data = 3'b111;
			92	: image_pixel_data = 3'b111;
			93	: image_pixel_data = 3'b111;
			94	: image_pixel_data = 3'b111;
			95	: image_pixel_data = 3'b111;
			96	: image_pixel_data = 3'b111;
			97	: image_pixel_data = 3'b111;
			98	: image_pixel_data = 3'b111;
			99	: image_pixel_data = 3'b111;
			100	: image_pixel_data = 3'b111;
			101	: image_pixel_data = 3'b000;
			102	: image_pixel_data = 3'b111;
			103	: image_pixel_data = 3'b111;
			104	: image_pixel_data = 3'b111;
			105	: image_pixel_data = 3'b111;
			106	: image_pixel_data = 3'b110;
			107	: image_pixel_data = 3'b110;
			108	: image_pixel_data = 3'b111;
			109	: image_pixel_data = 3'b111;
			110	: image_pixel_data = 3'b111;
			111	: image_pixel_data = 3'b111;
			112	: image_pixel_data = 3'b111;
			113	: image_pixel_data = 3'b111;
			114	: image_pixel_data = 3'b111;
			115	: image_pixel_data = 3'b111;
			116	: image_pixel_data = 3'b111;
			117	: image_pixel_data = 3'b000;
			118	: image_pixel_data = 3'b000;
			119	: image_pixel_data = 3'b000;
			120	: image_pixel_data = 3'b000;
			121	: image_pixel_data = 3'b111;
			122	: image_pixel_data = 3'b000;
			123	: image_pixel_data = 3'b111;
			124	: image_pixel_data = 3'b111;
			125	: image_pixel_data = 3'b111;
			126	: image_pixel_data = 3'b111;
			127	: image_pixel_data = 3'b111;
			128	: image_pixel_data = 3'b111;
			129	: image_pixel_data = 3'b111;
			130	: image_pixel_data = 3'b111;
			131	: image_pixel_data = 3'b111;
			132	: image_pixel_data = 3'b111;
			133	: image_pixel_data = 3'b111;
			134	: image_pixel_data = 3'b000;
			135	: image_pixel_data = 3'b000;
			136	: image_pixel_data = 3'b000;
			137	: image_pixel_data = 3'b111;
			138	: image_pixel_data = 3'b000;
			139	: image_pixel_data = 3'b111;
			140	: image_pixel_data = 3'b111;
			141	: image_pixel_data = 3'b111;
			142	: image_pixel_data = 3'b111;
			143	: image_pixel_data = 3'b111;
			144	: image_pixel_data = 3'b111;
			145	: image_pixel_data = 3'b111;
			146	: image_pixel_data = 3'b111;
			147	: image_pixel_data = 3'b111;
			148	: image_pixel_data = 3'b111;
			149	: image_pixel_data = 3'b111;
			150	: image_pixel_data = 3'b000;
			151	: image_pixel_data = 3'b000;
			152	: image_pixel_data = 3'b000;
			153	: image_pixel_data = 3'b111;
			154	: image_pixel_data = 3'b000;
			155	: image_pixel_data = 3'b111;
			156	: image_pixel_data = 3'b111;
			157	: image_pixel_data = 3'b111;
			158	: image_pixel_data = 3'b111;
			159	: image_pixel_data = 3'b111;
			160	: image_pixel_data = 3'b111;
			161	: image_pixel_data = 3'b111;
			162	: image_pixel_data = 3'b111;
			163	: image_pixel_data = 3'b111;
			164	: image_pixel_data = 3'b111;
			165	: image_pixel_data = 3'b111;
			166	: image_pixel_data = 3'b000;
			167	: image_pixel_data = 3'b111;
			168	: image_pixel_data = 3'b000;
			169	: image_pixel_data = 3'b111;
			170	: image_pixel_data = 3'b000;
			171	: image_pixel_data = 3'b111;
			172	: image_pixel_data = 3'b111;
			173	: image_pixel_data = 3'b111;
			174	: image_pixel_data = 3'b111;
			175	: image_pixel_data = 3'b111;
			176	: image_pixel_data = 3'b111;
			177	: image_pixel_data = 3'b111;
			178	: image_pixel_data = 3'b111;
			179	: image_pixel_data = 3'b111;
			180	: image_pixel_data = 3'b111;
			181	: image_pixel_data = 3'b111;
			182	: image_pixel_data = 3'b000;
			183	: image_pixel_data = 3'b111;
			184	: image_pixel_data = 3'b111;
			185	: image_pixel_data = 3'b111;
			186	: image_pixel_data = 3'b000;
			187	: image_pixel_data = 3'b111;
			188	: image_pixel_data = 3'b111;
			189	: image_pixel_data = 3'b111;
			190	: image_pixel_data = 3'b111;
			191	: image_pixel_data = 3'b111;
			192	: image_pixel_data = 3'b111;
			193	: image_pixel_data = 3'b111;
			194	: image_pixel_data = 3'b111;
			195	: image_pixel_data = 3'b111;
			196	: image_pixel_data = 3'b111;
			197	: image_pixel_data = 3'b111;
			198	: image_pixel_data = 3'b000;
			199	: image_pixel_data = 3'b000;
			200	: image_pixel_data = 3'b111;
			201	: image_pixel_data = 3'b111;
			202	: image_pixel_data = 3'b000;
			203	: image_pixel_data = 3'b111;
			204	: image_pixel_data = 3'b111;
			205	: image_pixel_data = 3'b111;
			206	: image_pixel_data = 3'b111;
			207	: image_pixel_data = 3'b111;
			208	: image_pixel_data = 3'b111;
			209	: image_pixel_data = 3'b111;
			210	: image_pixel_data = 3'b111;
			211	: image_pixel_data = 3'b111;
			212	: image_pixel_data = 3'b111;
			213	: image_pixel_data = 3'b111;
			214	: image_pixel_data = 3'b111;
			215	: image_pixel_data = 3'b000;
			216	: image_pixel_data = 3'b000;
			217	: image_pixel_data = 3'b000;
			218	: image_pixel_data = 3'b110;
			219	: image_pixel_data = 3'b110;
			220	: image_pixel_data = 3'b111;
			221	: image_pixel_data = 3'b111;
			222	: image_pixel_data = 3'b111;
			223	: image_pixel_data = 3'b111;
			224	: image_pixel_data = 3'b111;
			225	: image_pixel_data = 3'b111;
			226	: image_pixel_data = 3'b111;
			227	: image_pixel_data = 3'b111;
			228	: image_pixel_data = 3'b111;
			229	: image_pixel_data = 3'b111;
			230	: image_pixel_data = 3'b111;
			231	: image_pixel_data = 3'b111;
			232	: image_pixel_data = 3'b111;
			233	: image_pixel_data = 3'b111;
			234	: image_pixel_data = 3'b111;
			235	: image_pixel_data = 3'b111;
			236	: image_pixel_data = 3'b111;
			237	: image_pixel_data = 3'b111;
			238	: image_pixel_data = 3'b111;
			239	: image_pixel_data = 3'b111;
			240	: image_pixel_data = 3'b111;
			241	: image_pixel_data = 3'b111;
			242	: image_pixel_data = 3'b111;
			243	: image_pixel_data = 3'b111;
			244	: image_pixel_data = 3'b111;
			245	: image_pixel_data = 3'b111;
			246	: image_pixel_data = 3'b111;
			247	: image_pixel_data = 3'b111;
			248	: image_pixel_data = 3'b111;
			249	: image_pixel_data = 3'b111;
			250	: image_pixel_data = 3'b111;
			251	: image_pixel_data = 3'b111;
			252	: image_pixel_data = 3'b111;
			253	: image_pixel_data = 3'b111;
			254	: image_pixel_data = 3'b111;
			255	: image_pixel_data = 3'b111;
		endcase
	end
endtask

task image3_data;
	input [7:0] image_pixel_addr;
	output [2:0] image_pixel_data;
	reg [2:0] image_pixel_data;
	begin
		case (image_pixel_addr)
			0	: image_pixel_data = 3'b111;
			1	: image_pixel_data = 3'b111;
			2	: image_pixel_data = 3'b111;
			3	: image_pixel_data = 3'b111;
			4	: image_pixel_data = 3'b111;
			5	: image_pixel_data = 3'b111;
			6	: image_pixel_data = 3'b111;
			7	: image_pixel_data = 3'b111;
			8	: image_pixel_data = 3'b111;
			9	: image_pixel_data = 3'b111;
			10	: image_pixel_data = 3'b111;
			11	: image_pixel_data = 3'b111;
			12	: image_pixel_data = 3'b111;
			13	: image_pixel_data = 3'b111;
			14	: image_pixel_data = 3'b111;
			15	: image_pixel_data = 3'b111;
			16	: image_pixel_data = 3'b111;
			17	: image_pixel_data = 3'b111;
			18	: image_pixel_data = 3'b111;
			19	: image_pixel_data = 3'b111;
			20	: image_pixel_data = 3'b111;
			21	: image_pixel_data = 3'b111;
			22	: image_pixel_data = 3'b000;
			23	: image_pixel_data = 3'b000;
			24	: image_pixel_data = 3'b000;
			25	: image_pixel_data = 3'b000;
			26	: image_pixel_data = 3'b111;
			27	: image_pixel_data = 3'b111;
			28	: image_pixel_data = 3'b111;
			29	: image_pixel_data = 3'b111;
			30	: image_pixel_data = 3'b111;
			31	: image_pixel_data = 3'b111;
			32	: image_pixel_data = 3'b111;
			33	: image_pixel_data = 3'b111;
			34	: image_pixel_data = 3'b111;
			35	: image_pixel_data = 3'b111;
			36	: image_pixel_data = 3'b111;
			37	: image_pixel_data = 3'b000;
			38	: image_pixel_data = 3'b000;
			39	: image_pixel_data = 3'b000;
			40	: image_pixel_data = 3'b000;
			41	: image_pixel_data = 3'b000;
			42	: image_pixel_data = 3'b000;
			43	: image_pixel_data = 3'b111;
			44	: image_pixel_data = 3'b111;
			45	: image_pixel_data = 3'b111;
			46	: image_pixel_data = 3'b111;
			47	: image_pixel_data = 3'b111;
			48	: image_pixel_data = 3'b111;
			49	: image_pixel_data = 3'b111;
			50	: image_pixel_data = 3'b111;
			51	: image_pixel_data = 3'b111;
			52	: image_pixel_data = 3'b000;
			53	: image_pixel_data = 3'b000;
			54	: image_pixel_data = 3'b000;
			55	: image_pixel_data = 3'b000;
			56	: image_pixel_data = 3'b000;
			57	: image_pixel_data = 3'b000;
			58	: image_pixel_data = 3'b000;
			59	: image_pixel_data = 3'b000;
			60	: image_pixel_data = 3'b111;
			61	: image_pixel_data = 3'b111;
			62	: image_pixel_data = 3'b111;
			63	: image_pixel_data = 3'b111;
			64	: image_pixel_data = 3'b111;
			65	: image_pixel_data = 3'b111;
			66	: image_pixel_data = 3'b111;
			67	: image_pixel_data = 3'b111;
			68	: image_pixel_data = 3'b000;
			69	: image_pixel_data = 3'b000;
			70	: image_pixel_data = 3'b000;
			71	: image_pixel_data = 3'b000;
			72	: image_pixel_data = 3'b000;
			73	: image_pixel_data = 3'b000;
			74	: image_pixel_data = 3'b000;
			75	: image_pixel_data = 3'b000;
			76	: image_pixel_data = 3'b111;
			77	: image_pixel_data = 3'b111;
			78	: image_pixel_data = 3'b111;
			79	: image_pixel_data = 3'b111;
			80	: image_pixel_data = 3'b111;
			81	: image_pixel_data = 3'b111;
			82	: image_pixel_data = 3'b111;
			83	: image_pixel_data = 3'b111;
			84	: image_pixel_data = 3'b000;
			85	: image_pixel_data = 3'b000;
			86	: image_pixel_data = 3'b000;
			87	: image_pixel_data = 3'b000;
			88	: image_pixel_data = 3'b000;
			89	: image_pixel_data = 3'b000;
			90	: image_pixel_data = 3'b000;
			91	: image_pixel_data = 3'b000;
			92	: image_pixel_data = 3'b111;
			93	: image_pixel_data = 3'b111;
			94	: image_pixel_data = 3'b111;
			95	: image_pixel_data = 3'b111;
			96	: image_pixel_data = 3'b111;
			97	: image_pixel_data = 3'b111;
			98	: image_pixel_data = 3'b111;
			99	: image_pixel_data = 3'b000;
			100	: image_pixel_data = 3'b000;
			101	: image_pixel_data = 3'b000;
			102	: image_pixel_data = 3'b000;
			103	: image_pixel_data = 3'b000;
			104	: image_pixel_data = 3'b000;
			105	: image_pixel_data = 3'b000;
			106	: image_pixel_data = 3'b000;
			107	: image_pixel_data = 3'b000;
			108	: image_pixel_data = 3'b000;
			109	: image_pixel_data = 3'b111;
			110	: image_pixel_data = 3'b111;
			111	: image_pixel_data = 3'b111;
			112	: image_pixel_data = 3'b111;
			113	: image_pixel_data = 3'b111;
			114	: image_pixel_data = 3'b000;
			115	: image_pixel_data = 3'b000;
			116	: image_pixel_data = 3'b000;
			117	: image_pixel_data = 3'b000;
			118	: image_pixel_data = 3'b000;
			119	: image_pixel_data = 3'b000;
			120	: image_pixel_data = 3'b000;
			121	: image_pixel_data = 3'b000;
			122	: image_pixel_data = 3'b000;
			123	: image_pixel_data = 3'b000;
			124	: image_pixel_data = 3'b000;
			125	: image_pixel_data = 3'b000;
			126	: image_pixel_data = 3'b111;
			127	: image_pixel_data = 3'b111;
			128	: image_pixel_data = 3'b111;
			129	: image_pixel_data = 3'b111;
			130	: image_pixel_data = 3'b000;
			131	: image_pixel_data = 3'b000;
			132	: image_pixel_data = 3'b000;
			133	: image_pixel_data = 3'b000;
			134	: image_pixel_data = 3'b000;
			135	: image_pixel_data = 3'b000;
			136	: image_pixel_data = 3'b000;
			137	: image_pixel_data = 3'b000;
			138	: image_pixel_data = 3'b000;
			139	: image_pixel_data = 3'b000;
			140	: image_pixel_data = 3'b000;
			141	: image_pixel_data = 3'b000;
			142	: image_pixel_data = 3'b111;
			143	: image_pixel_data = 3'b111;
			144	: image_pixel_data = 3'b111;
			145	: image_pixel_data = 3'b111;
			146	: image_pixel_data = 3'b000;
			147	: image_pixel_data = 3'b111;
			148	: image_pixel_data = 3'b000;
			149	: image_pixel_data = 3'b000;
			150	: image_pixel_data = 3'b000;
			151	: image_pixel_data = 3'b000;
			152	: image_pixel_data = 3'b000;
			153	: image_pixel_data = 3'b000;
			154	: image_pixel_data = 3'b000;
			155	: image_pixel_data = 3'b000;
			156	: image_pixel_data = 3'b111;
			157	: image_pixel_data = 3'b000;
			158	: image_pixel_data = 3'b111;
			159	: image_pixel_data = 3'b111;
			160	: image_pixel_data = 3'b111;
			161	: image_pixel_data = 3'b111;
			162	: image_pixel_data = 3'b111;
			163	: image_pixel_data = 3'b111;
			164	: image_pixel_data = 3'b000;
			165	: image_pixel_data = 3'b000;
			166	: image_pixel_data = 3'b000;
			167	: image_pixel_data = 3'b000;
			168	: image_pixel_data = 3'b000;
			169	: image_pixel_data = 3'b000;
			170	: image_pixel_data = 3'b000;
			171	: image_pixel_data = 3'b000;
			172	: image_pixel_data = 3'b111;
			173	: image_pixel_data = 3'b111;
			174	: image_pixel_data = 3'b111;
			175	: image_pixel_data = 3'b111;
			176	: image_pixel_data = 3'b111;
			177	: image_pixel_data = 3'b111;
			178	: image_pixel_data = 3'b111;
			179	: image_pixel_data = 3'b111;
			180	: image_pixel_data = 3'b000;
			181	: image_pixel_data = 3'b000;
			182	: image_pixel_data = 3'b000;
			183	: image_pixel_data = 3'b000;
			184	: image_pixel_data = 3'b000;
			185	: image_pixel_data = 3'b000;
			186	: image_pixel_data = 3'b000;
			187	: image_pixel_data = 3'b000;
			188	: image_pixel_data = 3'b111;
			189	: image_pixel_data = 3'b111;
			190	: image_pixel_data = 3'b111;
			191	: image_pixel_data = 3'b111;
			192	: image_pixel_data = 3'b111;
			193	: image_pixel_data = 3'b111;
			194	: image_pixel_data = 3'b111;
			195	: image_pixel_data = 3'b111;
			196	: image_pixel_data = 3'b000;
			197	: image_pixel_data = 3'b000;
			198	: image_pixel_data = 3'b000;
			199	: image_pixel_data = 3'b000;
			200	: image_pixel_data = 3'b000;
			201	: image_pixel_data = 3'b000;
			202	: image_pixel_data = 3'b000;
			203	: image_pixel_data = 3'b000;
			204	: image_pixel_data = 3'b111;
			205	: image_pixel_data = 3'b111;
			206	: image_pixel_data = 3'b111;
			207	: image_pixel_data = 3'b111;
			208	: image_pixel_data = 3'b111;
			209	: image_pixel_data = 3'b111;
			210	: image_pixel_data = 3'b111;
			211	: image_pixel_data = 3'b111;
			212	: image_pixel_data = 3'b111;
			213	: image_pixel_data = 3'b110;
			214	: image_pixel_data = 3'b110;
			215	: image_pixel_data = 3'b000;
			216	: image_pixel_data = 3'b000;
			217	: image_pixel_data = 3'b110;
			218	: image_pixel_data = 3'b110;
			219	: image_pixel_data = 3'b111;
			220	: image_pixel_data = 3'b111;
			221	: image_pixel_data = 3'b111;
			222	: image_pixel_data = 3'b111;
			223	: image_pixel_data = 3'b111;
			224	: image_pixel_data = 3'b111;
			225	: image_pixel_data = 3'b111;
			226	: image_pixel_data = 3'b111;
			227	: image_pixel_data = 3'b111;
			228	: image_pixel_data = 3'b111;
			229	: image_pixel_data = 3'b111;
			230	: image_pixel_data = 3'b111;
			231	: image_pixel_data = 3'b111;
			232	: image_pixel_data = 3'b111;
			233	: image_pixel_data = 3'b111;
			234	: image_pixel_data = 3'b111;
			235	: image_pixel_data = 3'b111;
			236	: image_pixel_data = 3'b111;
			237	: image_pixel_data = 3'b111;
			238	: image_pixel_data = 3'b111;
			239	: image_pixel_data = 3'b111;
			240	: image_pixel_data = 3'b111;
			241	: image_pixel_data = 3'b111;
			242	: image_pixel_data = 3'b111;
			243	: image_pixel_data = 3'b111;
			244	: image_pixel_data = 3'b111;
			245	: image_pixel_data = 3'b111;
			246	: image_pixel_data = 3'b111;
			247	: image_pixel_data = 3'b111;
			248	: image_pixel_data = 3'b111;
			249	: image_pixel_data = 3'b111;
			250	: image_pixel_data = 3'b111;
			251	: image_pixel_data = 3'b111;
			252	: image_pixel_data = 3'b111;
			253	: image_pixel_data = 3'b111;
			254	: image_pixel_data = 3'b111;
			255	: image_pixel_data = 3'b111;
		endcase
	end
endtask

always @(*) begin
	//Sync the current image.
	current_image = image_index;
	//Get the image index.
	case (current_image)
		// Image #0
		0: begin
			image0_data(func2_pixel_addr, func2_pixel_data);
			image0_data(func3_pixel_addr, func3_pixel_data);
		end
		// Image #1
		1: begin
			image1_data(func2_pixel_addr, func2_pixel_data);
			image1_data(func3_pixel_addr, func3_pixel_data);
		end
		// Image #2
		2: begin
			image2_data(func2_pixel_addr, func2_pixel_data);
			image2_data(func3_pixel_addr, func3_pixel_data);
		end
		// Image #4
		3: begin
			image3_data(func2_pixel_addr, func2_pixel_data);
			image3_data(func3_pixel_addr, func3_pixel_data);
		end
	endcase
end

endmodule